input component

component()
